package Instance_Incoherent where

import IncoherentBase
import Vector

class incoherent DependingIncoherent a where
  dependMethod :: a -> String

instance (IncoherentBase a) => DependingIncoherent a where
  dependMethod x = "incoherent " +++ printType (typeOf x) +++ ": " +++ baseMethod x

testByteDirect :: String
testByteDirect =
  let v :: Vector 4 Byte
      v = replicate 0
  in dependMethod v

testIntDirect :: String
testIntDirect =
  let v :: Vector 4 (Int 8)
      v = replicate 0
  in dependMethod v

useGeneric :: Vector n a -> String
useGeneric v = dependMethod v

testByteViaGeneric :: String
testByteViaGeneric = useGeneric ((replicate 0) :: Vector 4 Byte)

sysInstance_Incoherent :: Module Empty
sysInstance_Incoherent = module
  rules
    "show": when True ==> do
      $display "Byte direct: " testByteDirect
      $display "Int direct: " testIntDirect
      $display "Byte via generic: " testByteViaGeneric
      $finish 0
